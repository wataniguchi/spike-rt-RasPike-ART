/*
 *  TOPPERS Software
 *      Toyohashi Open Platform for Embedded Real-Time Systems
 *
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015-2022 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 *
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 *
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 */

/*
 *    シリアルインタフェースドライバのコンポーネント記述ファイル
 */

/*
 *  シリアルインタフェースドライバをTECSを用いずに呼び出すためにも必要
 *  な定義の取込み
 */
import_C("syssvc/serial.h");

/*
 *  シリアルインタフェースドライバのターゲット依存部が提供する関数
 */
signature sSIOAsyncPort {
  void  open(void);
  void  close(void);
  void  putNotify(void);
  void  enableCBR([in] uint_t cbrtn);
  void  disableCBR([in] uint_t cbrtn);
};

/*
 *  コールバックルーチンの識別番号（cbrtnパラメータに用いる）
 */
const uint_t SIOAsyncSendPop = 1;   /* 送信可能コールバック */
const uint_t SIOAsyncReceivePush = 2; /* 受信通知コールバック */

/*
 *  ターゲット依存部からのコールバック
 */
[callback]
signature sSIOAsyncCBR {
  ER_UINT popSend([out] char *dst);
  //ER_UINT popSend([out] char *dst_data, [in] uint_t max_size);
  ER_UINT pushReceive([in] char src);
  //ER_UINT pushReceive([in] const char *src_data, [in] uint_t size);
  ER_UINT sizeSend(void);
};

/*
 *  シリアルポートの制御部のセルタイプ
 */
celltype tSerialAsyncPortMain {
  entry sSerialPort     eSerialPort;
  entry snSerialPortManage  enSerialPortManage;

  call  sSIOAsyncPort cSIOPort;     /* 簡易SIOドライバとの接続 */
  entry sSIOAsyncCBR  eSIOCBR;

  call  sSemaphore  cSendSemaphore;   /* 送信用セマフォとの接続 */
  call  sSemaphore  cReceiveSemaphore;  /* 受信用セマフォとの接続 */

  attr {
    uint_t  receiveBufferSize = 256;  /* 受信バッファサイズ */
    uint_t  sendBufferSize = 256;   /* 送信バッファサイズ */
  };
  var {
    bool_t  openFlag = C_EXP("false");  /* オープン済みフラグ */
    bool_t  errorFlag;          /* エラーフラグ */
    uint_t  ioControl;          /* 動作制御の設定値 */

    [size_is(receiveBufferSize)] char *receiveBuffer; /* 受信バッファ */
    uint_t  receiveReadPointer;     /* 受信バッファ読出しポインタ */
    uint_t  receiveWritePointer;    /* 受信バッファ書込みポインタ */
    uint_t  receiveCount;       /* 受信バッファ中の文字数 */

    [size_is(sendBufferSize)] char *sendBuffer;   /* 送信バッファ */
    uint_t  sendReadPointer;      /* 送信バッファ読出しポインタ */
    uint_t  sendWritePointer;     /* 送信バッファ書込みポインタ */
    uint_t  sendCount;          /* 送信バッファ中の文字数 */
  };
};

/*
 *  シリアルポートドライバ（複合セル）のセルタイプ
 *
 *  シリアルポートの制御部と，それが使用する2つのセマフォ（受信用と送
 *  信用）を複合化して，1つのコンポーネントとしている．
 */
composite tSerialAsyncPort {
  entry sSerialPort     eSerialPort;
  entry snSerialPortManage  enSerialPortManage;

  call  sSIOAsyncPort   cSIOPort;   /* 簡易SIOドライバとの接続 */
  entry sSIOAsyncCBR    eSIOCBR;

  attr {
    uint_t  receiveBufferSize = 256;  /* 受信バッファサイズ */
    uint_t  sendBufferSize = 256;   /* 送信バッファサイズ */
  };

  /* 受信用のセマフォ */
  cell tSemaphore ReceiveSemaphore {
    attribute = C_EXP("TA_NULL");
    initialCount = 0;
    maxCount =1;
  };

  /* 送信用のセマフォ */
  cell tSemaphore SendSemaphore {
    attribute = C_EXP("TA_NULL");
    initialCount = 1;
    maxCount =1;
  };

  /* シリアルポートの制御部 */
  cell tSerialAsyncPortMain SerialPortMain {
    /* セマフォとの結合 */
    cReceiveSemaphore  = ReceiveSemaphore.eSemaphore;
    cSendSemaphore     = SendSemaphore.eSemaphore;

    /* 呼び口のエクスポート */
    cSIOPort          => composite.cSIOPort;

    /* 属性の継承 */
    receiveBufferSize = composite.receiveBufferSize;
    sendBufferSize    = composite.sendBufferSize;
  };

  /* 受け口のエクスポート */
  composite.eSerialPort        => SerialPortMain.eSerialPort;
  composite.enSerialPortManage => SerialPortMain.enSerialPortManage;
  composite.eSIOCBR            => SerialPortMain.eSIOCBR;
};
